package Rng;

import GetPut::*;
import FIFOF::*;
import LFSR::*;
import FixedPoint::*;
import Vector::*;


module mkSqrtPipeline#(numeric n) ();

endmodule

(* synthesize *)
module mkGaussianRNG ();

endmodule

endpackage