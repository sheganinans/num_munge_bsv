package LnPipeline;

import FixedPoint::*;
import FIFOF::*;

`include "DEFNS.defines"

typedef FixedPoint#(`FixPointSizes) FXP;

endpackage
